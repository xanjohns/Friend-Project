 logic test;
           logic clk;
  
  
logic clk2;
   logic newtest;
