 logic test;
           logic clk;


logic clk2;
