 logic test;

   logic test2;
            logic test4;
